module MIPS()
reg MuxCtrl;

initial
begin
MuxCtrl<=0;
end
endmodule
